

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity main2 is
port();
end main2;

architecture Behavioral of main2 is
begin

end Behavioral;


